module circuit_a(
    // Declare inputs
    // Declare Y output
    //test
);

    // Enter logic equation here

endmodule
